../../../hdl/wb_cdc/wb_cdc.vhd